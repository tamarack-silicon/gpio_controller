module gpio_controller_verif_tb;

	initial begin
		uvm_pkg::run_test();
	end

endmodule // gpio_controller_verif_tb
