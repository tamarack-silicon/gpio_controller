module gpio_controller;

endmodule // gpio_controller
