module gpio_controller_tb;

endmodule // gpio_controller_tb
